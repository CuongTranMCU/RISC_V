module Adder(In1,In2,Out);
output [31:0] Out;
input [31:0] In1,In2;
assign Out = In1 + In2;
endmodule
